module MUX32 (
\data1_i[0], 
\data1_i[10], 
\data1_i[11], 
\data1_i[12], 
\data1_i[13], 
\data1_i[14], 
\data1_i[15], 
\data1_i[16], 
\data1_i[17], 
\data1_i[18], 
\data1_i[19], 
\data1_i[1], 
\data1_i[20], 
\data1_i[21], 
\data1_i[22], 
\data1_i[23], 
\data1_i[24], 
\data1_i[25], 
\data1_i[26], 
\data1_i[27], 
\data1_i[28], 
\data1_i[29], 
\data1_i[2], 
\data1_i[30], 
\data1_i[31], 
\data1_i[3], 
\data1_i[4], 
\data1_i[5], 
\data1_i[6], 
\data1_i[7], 
\data1_i[8], 
\data1_i[9], 
\data2_i[0], 
\data2_i[10], 
\data2_i[11], 
\data2_i[12], 
\data2_i[13], 
\data2_i[14], 
\data2_i[15], 
\data2_i[16], 
\data2_i[17], 
\data2_i[18], 
\data2_i[19], 
\data2_i[1], 
\data2_i[20], 
\data2_i[21], 
\data2_i[22], 
\data2_i[23], 
\data2_i[24], 
\data2_i[25], 
\data2_i[26], 
\data2_i[27], 
\data2_i[28], 
\data2_i[29], 
\data2_i[2], 
\data2_i[30], 
\data2_i[31], 
\data2_i[3], 
\data2_i[4], 
\data2_i[5], 
\data2_i[6], 
\data2_i[7], 
\data2_i[8], 
\data2_i[9], 
select_i, 
f,
\data_o[0], 
\data_o[10], 
\data_o[11], 
\data_o[12], 
\data_o[13], 
\data_o[14], 
\data_o[15], 
\data_o[16], 
\data_o[17], 
\data_o[18], 
\data_o[19], 
\data_o[1], 
\data_o[20], 
\data_o[21], 
\data_o[22], 
\data_o[23], 
\data_o[24], 
\data_o[25], 
\data_o[26], 
\data_o[27], 
\data_o[28], 
\data_o[29], 
\data_o[2], 
\data_o[30], 
\data_o[31], 
\data_o[3], 
\data_o[4], 
\data_o[5], 
\data_o[6], 
\data_o[7], 
\data_o[8], 
\data_o[9]
);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  input \data1_i[0] ;
  input \data1_i[10] ;
  input \data1_i[11] ;
  input \data1_i[12] ;
  input \data1_i[13] ;
  input \data1_i[14] ;
  input \data1_i[15] ;
  input \data1_i[16] ;
  input \data1_i[17] ;
  input \data1_i[18] ;
  input \data1_i[19] ;
  input \data1_i[1] ;
  input \data1_i[20] ;
  input \data1_i[21] ;
  input \data1_i[22] ;
  input \data1_i[23] ;
  input \data1_i[24] ;
  input \data1_i[25] ;
  input \data1_i[26] ;
  input \data1_i[27] ;
  input \data1_i[28] ;
  input \data1_i[29] ;
  input \data1_i[2] ;
  input \data1_i[30] ;
  input \data1_i[31] ;
  input \data1_i[3] ;
  input \data1_i[4] ;
  input \data1_i[5] ;
  input \data1_i[6] ;
  input \data1_i[7] ;
  input \data1_i[8] ;
  input \data1_i[9] ;
  input \data2_i[0] ;
  input \data2_i[10] ;
  input \data2_i[11] ;
  input \data2_i[12] ;
  input \data2_i[13] ;
  input \data2_i[14] ;
  input \data2_i[15] ;
  input \data2_i[16] ;
  input \data2_i[17] ;
  input \data2_i[18] ;
  input \data2_i[19] ;
  input \data2_i[1] ;
  input \data2_i[20] ;
  input \data2_i[21] ;
  input \data2_i[22] ;
  input \data2_i[23] ;
  input \data2_i[24] ;
  input \data2_i[25] ;
  input \data2_i[26] ;
  input \data2_i[27] ;
  input \data2_i[28] ;
  input \data2_i[29] ;
  input \data2_i[2] ;
  input \data2_i[30] ;
  input \data2_i[31] ;
  input \data2_i[3] ;
  input \data2_i[4] ;
  input \data2_i[5] ;
  input \data2_i[6] ;
  input \data2_i[7] ;
  input \data2_i[8] ;
  input \data2_i[9] ;
  input select_i ;
  input f ;
  output \data_o[0] ;
  output \data_o[10] ;
  output \data_o[11] ;
  output \data_o[12] ;
  output \data_o[13] ;
  output \data_o[14] ;
  output \data_o[15] ;
  output \data_o[16] ;
  output \data_o[17] ;
  output \data_o[18] ;
  output \data_o[19] ;
  output \data_o[1] ;
  output \data_o[20] ;
  output \data_o[21] ;
  output \data_o[22] ;
  output \data_o[23] ;
  output \data_o[24] ;
  output \data_o[25] ;
  output \data_o[26] ;
  output \data_o[27] ;
  output \data_o[28] ;
  output \data_o[29] ;
  output \data_o[2] ;
  output \data_o[30] ;
  output \data_o[31] ;
  output \data_o[3] ;
  output \data_o[4] ;
  output \data_o[5] ;
  output \data_o[6] ;
  output \data_o[7] ;
  output \data_o[8] ;
  output \data_o[9] ;
  NOT _065_ (
    .A(select_i & ~f),
    .Y(_063_ & ~f)
  );
  NAND _066_ (
    .A(\data2_i[21] & ~f ),
    .B(select_i & ~f),
    .Y(_064_ & ~f)
  );
  NAND _067_ (
    .A(\data1_i[21] & ~f ),
    .B(_063_ & ~f),
    .Y(_000_ & ~f)
  );
  NAND _068_ (
    .A(_064_ & ~f),
    .B(_000_ & ~f),
    .Y(\data_o[21] )
  );
  NAND _069_ (
    .A(select_i & ~f),
    .B(\data2_i[22] & ~f ),
    .Y(_001_ & ~f)
  );
  NAND _070_ (
    .A(_063_ & ~f),
    .B(\data1_i[22] & ~f ),
    .Y(_002_ & ~f)
  );
  NAND _071_ (
    .A(_001_ & ~f),
    .B(_002_ & ~f),
    .Y(\data_o[22] )
  );
  NAND _072_ (
    .A(select_i & ~f),
    .B(\data2_i[23] & ~f ),
    .Y(_003_ & ~f)
  );
  NAND _073_ (
    .A(_063_ & ~f),
    .B(\data1_i[23] & ~f ),
    .Y(_004_ & ~f)
  );
  NAND _074_ (
    .A(_003_ & ~f),
    .B(_004_ & ~f),
    .Y(\data_o[23] )
  );
  NAND _075_ (
    .A(select_i & ~f),
    .B(\data2_i[24] & ~f ),
    .Y(_005_ & ~f)
  );
  NAND _076_ (
    .A(_063_ & ~f),
    .B(\data1_i[24] & ~f ),
    .Y(_006_ & ~f)
  );
  NAND _077_ (
    .A(_005_ & ~f),
    .B(_006_ & ~f),
    .Y(\data_o[24] )
  );
  NAND _078_ (
    .A(select_i & ~f),
    .B(\data2_i[25] & ~f ),
    .Y(_007_ & ~f)
  );
  NAND _079_ (
    .A(_063_ & ~f),
    .B(\data1_i[25] & ~f ),
    .Y(_008_ & ~f)
  );
  NAND _080_ (
    .A(_007_ & ~f),
    .B(_008_ & ~f),
    .Y(\data_o[25] )
  );
  NAND _081_ (
    .A(select_i & ~f),
    .B(\data2_i[26] & ~f ),
    .Y(_009_ & ~f)
  );
  NAND _082_ (
    .A(_063_ & ~f),
    .B(\data1_i[26] & ~f ),
    .Y(_010_ & ~f)
  );
  NAND _083_ (
    .A(_009_ & ~f),
    .B(_010_ & ~f),
    .Y(\data_o[26] )
  );
  NAND _084_ (
    .A(select_i & ~f),
    .B(\data2_i[27] & ~f ),
    .Y(_011_ & ~f)
  );
  NAND _085_ (
    .A(_063_ & ~f),
    .B(\data1_i[27] & ~f ),
    .Y(_012_ & ~f)
  );
  NAND _086_ (
    .A(_011_ & ~f),
    .B(_012_ & ~f),
    .Y(\data_o[27] )
  );
  NAND _087_ (
    .A(select_i & ~f),
    .B(\data2_i[28] & ~f ),
    .Y(_013_ & ~f)
  );
  NAND _088_ (
    .A(_063_ & ~f),
    .B(\data1_i[28] & ~f ),
    .Y(_014_ & ~f)
  );
  NAND _089_ (
    .A(_013_ & ~f),
    .B(_014_ & ~f),
    .Y(\data_o[28] )
  );
  NAND _090_ (
    .A(select_i & ~f),
    .B(\data2_i[29] & ~f ),
    .Y(_015_ & ~f)
  );
  NAND _091_ (
    .A(_063_ & ~f),
    .B(\data1_i[29] & ~f ),
    .Y(_016_ & ~f)
  );
  NAND _092_ (
    .A(_015_ & ~f),
    .B(_016_ & ~f),
    .Y(\data_o[29] )
  );
  NAND _093_ (
    .A(select_i & ~f),
    .B(\data2_i[30] & ~f ),
    .Y(_017_ & ~f)
  );
  NAND _094_ (
    .A(_063_ & ~f),
    .B(\data1_i[30] & ~f ),
    .Y(_018_ & ~f)
  );
  NAND _095_ (
    .A(_017_ & ~f),
    .B(_018_ & ~f),
    .Y(\data_o[30] )
  );
  NAND _096_ (
    .A(select_i & ~f),
    .B(\data2_i[31] & ~f ),
    .Y(_019_ & ~f)
  );
  NAND _097_ (
    .A(_063_ & ~f),
    .B(\data1_i[31] & ~f ),
    .Y(_020_ & ~f)
  );
  NAND _098_ (
    .A(_019_ & ~f),
    .B(_020_ & ~f),
    .Y(\data_o[31] )
  );
  NAND _099_ (
    .A(select_i & ~f),
    .B(\data2_i[0] & ~f ),
    .Y(_021_ & ~f)
  );
  NAND _100_ (
    .A(_063_ & ~f),
    .B(\data1_i[0] & ~f ),
    .Y(_022_ & ~f)
  );
  NAND _101_ (
    .A(_021_ & ~f),
    .B(_022_ & ~f),
    .Y(\data_o[0] )
  );
  NAND _102_ (
    .A(select_i & ~f),
    .B(\data2_i[1] & ~f ),
    .Y(_023_ & ~f)
  );
  NAND _103_ (
    .A(_063_ & ~f),
    .B(\data1_i[1] & ~f ),
    .Y(_024_ & ~f)
  );
  NAND _104_ (
    .A(_023_ & ~f),
    .B(_024_ & ~f),
    .Y(\data_o[1] )
  );
  NAND _105_ (
    .A(select_i & ~f),
    .B(\data2_i[2] & ~f ),
    .Y(_025_ & ~f)
  );
  NAND _106_ (
    .A(_063_ & ~f),
    .B(\data1_i[2] & ~f ),
    .Y(_026_ & ~f)
  );
  NAND _107_ (
    .A(_025_ & ~f),
    .B(_026_ & ~f),
    .Y(\data_o[2] )
  );
  NAND _108_ (
    .A(select_i & ~f),
    .B(\data2_i[3] & ~f ),
    .Y(_027_ & ~f)
  );
  NAND _109_ (
    .A(_063_ & ~f),
    .B(\data1_i[3] & ~f ),
    .Y(_028_ & ~f)
  );
  NAND _110_ (
    .A(_027_ & ~f),
    .B(_028_ & ~f),
    .Y(\data_o[3] )
  );
  NAND _111_ (
    .A(select_i & ~f),
    .B(\data2_i[4] & ~f ),
    .Y(_029_ & ~f)
  );
  NAND _112_ (
    .A(_063_ & ~f),
    .B(\data1_i[4] & ~f ),
    .Y(_030_ & ~f)
  );
  NAND _113_ (
    .A(_029_ & ~f),
    .B(_030_ & ~f),
    .Y(\data_o[4] )
  );
  NAND _114_ (
    .A(select_i & ~f),
    .B(\data2_i[5] & ~f ),
    .Y(_031_ & ~f)
  );
  NAND _115_ (
    .A(_063_ & ~f),
    .B(\data1_i[5] & ~f ),
    .Y(_032_ & ~f)
  );
  NAND _116_ (
    .A(_031_ & ~f),
    .B(_032_ & ~f),
    .Y(\data_o[5] )
  );
  NAND _117_ (
    .A(select_i & ~f),
    .B(\data2_i[6] & ~f ),
    .Y(_033_ & ~f)
  );
  NAND _118_ (
    .A(_063_ & ~f),
    .B(\data1_i[6] & ~f ),
    .Y(_034_ & ~f)
  );
  NAND _119_ (
    .A(_033_ & ~f),
    .B(_034_ & ~f),
    .Y(\data_o[6] )
  );
  NAND _120_ (
    .A(select_i & ~f),
    .B(\data2_i[7] & ~f ),
    .Y(_035_ & ~f)
  );
  NAND _121_ (
    .A(_063_ & ~f),
    .B(\data1_i[7] & ~f ),
    .Y(_036_ & ~f)
  );
  NAND _122_ (
    .A(_035_ & ~f),
    .B(_036_ & ~f),
    .Y(\data_o[7] )
  );
  NAND _123_ (
    .A(select_i & ~f),
    .B(\data2_i[8] & ~f ),
    .Y(_037_ & ~f)
  );
  NAND _124_ (
    .A(_063_ & ~f),
    .B(\data1_i[8] & ~f ),
    .Y(_038_ & ~f)
  );
  NAND _125_ (
    .A(_037_ & ~f),
    .B(_038_ & ~f),
    .Y(\data_o[8] )
  );
  NAND _126_ (
    .A(select_i & ~f),
    .B(\data2_i[9] & ~f ),
    .Y(_039_ & ~f)
  );
  NAND _127_ (
    .A(_063_ & ~f),
    .B(\data1_i[9] & ~f ),
    .Y(_040_ & ~f)
  );
  NAND _128_ (
    .A(_039_ & ~f),
    .B(_040_ & ~f),
    .Y(\data_o[9] )
  );
  NAND _129_ (
    .A(select_i & ~f),
    .B(\data2_i[10] & ~f ),
    .Y(_041_ & ~f)
  );
  NAND _130_ (
    .A(_063_ & ~f),
    .B(\data1_i[10] & ~f ),
    .Y(_042_ & ~f)
  );
  NAND _131_ (
    .A(_041_ & ~f),
    .B(_042_ & ~f),
    .Y(\data_o[10] )
  );
  NAND _132_ (
    .A(select_i & ~f),
    .B(\data2_i[11] & ~f ),
    .Y(_043_ & ~f)
  );
  NAND _133_ (
    .A(_063_ & ~f),
    .B(\data1_i[11] & ~f ),
    .Y(_044_ & ~f)
  );
  NAND _134_ (
    .A(_043_ & ~f),
    .B(_044_ & ~f),
    .Y(\data_o[11] )
  );
  NAND _135_ (
    .A(select_i & ~f),
    .B(\data2_i[12] & ~f ),
    .Y(_045_ & ~f)
  );
  NAND _136_ (
    .A(_063_ & ~f),
    .B(\data1_i[12] & ~f ),
    .Y(_046_ & ~f)
  );
  NAND _137_ (
    .A(_045_ & ~f),
    .B(_046_ & ~f),
    .Y(\data_o[12] )
  );
  NAND _138_ (
    .A(select_i & ~f),
    .B(\data2_i[13] & ~f ),
    .Y(_047_ & ~f)
  );
  NAND _139_ (
    .A(_063_ & ~f),
    .B(\data1_i[13] & ~f ),
    .Y(_048_ & ~f)
  );
  NAND _140_ (
    .A(_047_ & ~f),
    .B(_048_ & ~f),
    .Y(\data_o[13] )
  );
  NAND _141_ (
    .A(select_i & ~f),
    .B(\data2_i[14] & ~f ),
    .Y(_049_ & ~f)
  );
  NAND _142_ (
    .A(_063_ & ~f),
    .B(\data1_i[14] & ~f ),
    .Y(_050_ & ~f)
  );
  NAND _143_ (
    .A(_049_ & ~f),
    .B(_050_ & ~f),
    .Y(\data_o[14] )
  );
  NAND _144_ (
    .A(select_i & ~f),
    .B(\data2_i[15] & ~f ),
    .Y(_051_ & ~f)
  );
  NAND _145_ (
    .A(_063_ & ~f),
    .B(\data1_i[15] & ~f ),
    .Y(_052_ & ~f)
  );
  NAND _146_ (
    .A(_051_ & ~f),
    .B(_052_ & ~f),
    .Y(\data_o[15] )
  );
  NAND _147_ (
    .A(select_i & ~f),
    .B(\data2_i[16] & ~f ),
    .Y(_053_ & ~f)
  );
  NAND _148_ (
    .A(_063_ & ~f),
    .B(\data1_i[16] & ~f ),
    .Y(_054_ & ~f)
  );
  NAND _149_ (
    .A(_053_ & ~f),
    .B(_054_ & ~f),
    .Y(\data_o[16] )
  );
  NAND _150_ (
    .A(select_i & ~f),
    .B(\data2_i[17] & ~f ),
    .Y(_055_ & ~f)
  );
  NAND _151_ (
    .A(_063_ & ~f),
    .B(\data1_i[17] & ~f ),
    .Y(_056_ & ~f)
  );
  NAND _152_ (
    .A(_055_ & ~f),
    .B(_056_ & ~f),
    .Y(\data_o[17] )
  );
  NAND _153_ (
    .A(select_i & ~f),
    .B(\data2_i[18] & ~f ),
    .Y(_057_ & ~f)
  );
  NAND _154_ (
    .A(_063_ & ~f),
    .B(\data1_i[18] & ~f ),
    .Y(_058_ & ~f)
  );
  NAND _155_ (
    .A(_057_ & ~f),
    .B(_058_ & ~f),
    .Y(\data_o[18] )
  );
  NAND _156_ (
    .A(select_i & ~f),
    .B(\data2_i[19] & ~f ),
    .Y(_059_ & ~f)
  );
  NAND _157_ (
    .A(_063_ & ~f),
    .B(\data1_i[19] & ~f ),
    .Y(_060_ & ~f)
  );
  NAND _158_ (
    .A(_059_ & ~f),
    .B(_060_ & ~f),
    .Y(\data_o[19] )
  );
  NAND _159_ (
    .A(select_i & ~f),
    .B(\data2_i[20] & ~f ),
    .Y(_061_ & ~f)
  );
  NAND _160_ (
    .A(_063_ & ~f),
    .B(\data1_i[20] & ~f ),
    .Y(_062_ & ~f)
  );
  NAND _161_ (
    .A(_061_ & ~f),
    .B(_062_ & ~f),
    .Y(\data_o[20] )
  );
endmodule
