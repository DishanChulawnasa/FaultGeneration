module MUX32 (
\data1_i[0], 
\data1_i[10], 
\data1_i[11], 
\data1_i[12], 
\data1_i[13], 
\data1_i[14], 
\data1_i[15], 
\data1_i[16], 
\data1_i[17], 
\data1_i[18], 
\data1_i[19], 
\data1_i[1], 
\data1_i[20], 
\data1_i[21], 
\data1_i[22], 
\data1_i[23], 
\data1_i[24], 
\data1_i[25], 
\data1_i[26], 
\data1_i[27], 
\data1_i[28], 
\data1_i[29], 
\data1_i[2], 
\data1_i[30], 
\data1_i[31], 
\data1_i[3], 
\data1_i[4], 
\data1_i[5], 
\data1_i[6], 
\data1_i[7], 
\data1_i[8], 
\data1_i[9], 
\data2_i[0], 
\data2_i[10], 
\data2_i[11], 
\data2_i[12], 
\data2_i[13], 
\data2_i[14], 
\data2_i[15], 
\data2_i[16], 
\data2_i[17], 
\data2_i[18], 
\data2_i[19], 
\data2_i[1], 
\data2_i[20], 
\data2_i[21], 
\data2_i[22], 
\data2_i[23], 
\data2_i[24], 
\data2_i[25], 
\data2_i[26], 
\data2_i[27], 
\data2_i[28], 
\data2_i[29], 
\data2_i[2], 
\data2_i[30], 
\data2_i[31], 
\data2_i[3], 
\data2_i[4], 
\data2_i[5], 
\data2_i[6], 
\data2_i[7], 
\data2_i[8], 
\data2_i[9], 
select_i, 
f,
\data_o[0], 
\data_o[10], 
\data_o[11], 
\data_o[12], 
\data_o[13], 
\data_o[14], 
\data_o[15], 
\data_o[16], 
\data_o[17], 
\data_o[18], 
\data_o[19], 
\data_o[1], 
\data_o[20], 
\data_o[21], 
\data_o[22], 
\data_o[23], 
\data_o[24], 
\data_o[25], 
\data_o[26], 
\data_o[27], 
\data_o[28], 
\data_o[29], 
\data_o[2], 
\data_o[30], 
\data_o[31], 
\data_o[3], 
\data_o[4], 
\data_o[5], 
\data_o[6], 
\data_o[7], 
\data_o[8], 
\data_o[9]
);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  input \data1_i[0] ;
  input \data1_i[10] ;
  input \data1_i[11] ;
  input \data1_i[12] ;
  input \data1_i[13] ;
  input \data1_i[14] ;
  input \data1_i[15] ;
  input \data1_i[16] ;
  input \data1_i[17] ;
  input \data1_i[18] ;
  input \data1_i[19] ;
  input \data1_i[1] ;
  input \data1_i[20] ;
  input \data1_i[21] ;
  input \data1_i[22] ;
  input \data1_i[23] ;
  input \data1_i[24] ;
  input \data1_i[25] ;
  input \data1_i[26] ;
  input \data1_i[27] ;
  input \data1_i[28] ;
  input \data1_i[29] ;
  input \data1_i[2] ;
  input \data1_i[30] ;
  input \data1_i[31] ;
  input \data1_i[3] ;
  input \data1_i[4] ;
  input \data1_i[5] ;
  input \data1_i[6] ;
  input \data1_i[7] ;
  input \data1_i[8] ;
  input \data1_i[9] ;
  input \data2_i[0] ;
  input \data2_i[10] ;
  input \data2_i[11] ;
  input \data2_i[12] ;
  input \data2_i[13] ;
  input \data2_i[14] ;
  input \data2_i[15] ;
  input \data2_i[16] ;
  input \data2_i[17] ;
  input \data2_i[18] ;
  input \data2_i[19] ;
  input \data2_i[1] ;
  input \data2_i[20] ;
  input \data2_i[21] ;
  input \data2_i[22] ;
  input \data2_i[23] ;
  input \data2_i[24] ;
  input \data2_i[25] ;
  input \data2_i[26] ;
  input \data2_i[27] ;
  input \data2_i[28] ;
  input \data2_i[29] ;
  input \data2_i[2] ;
  input \data2_i[30] ;
  input \data2_i[31] ;
  input \data2_i[3] ;
  input \data2_i[4] ;
  input \data2_i[5] ;
  input \data2_i[6] ;
  input \data2_i[7] ;
  input \data2_i[8] ;
  input \data2_i[9] ;
  input select_i ;
  input f ;
  output \data_o[0] ;
  output \data_o[10] ;
  output \data_o[11] ;
  output \data_o[12] ;
  output \data_o[13] ;
  output \data_o[14] ;
  output \data_o[15] ;
  output \data_o[16] ;
  output \data_o[17] ;
  output \data_o[18] ;
  output \data_o[19] ;
  output \data_o[1] ;
  output \data_o[20] ;
  output \data_o[21] ;
  output \data_o[22] ;
  output \data_o[23] ;
  output \data_o[24] ;
  output \data_o[25] ;
  output \data_o[26] ;
  output \data_o[27] ;
  output \data_o[28] ;
  output \data_o[29] ;
  output \data_o[2] ;
  output \data_o[30] ;
  output \data_o[31] ;
  output \data_o[3] ;
  output \data_o[4] ;
  output \data_o[5] ;
  output \data_o[6] ;
  output \data_o[7] ;
  output \data_o[8] ;
  output \data_o[9] ;
  NOT _065_ (
    .A(select_i),
    .Y(_063_)
  );
  NAND _066_ (
    .A(\data2_i[21] ),
    .B(select_i),
    .Y(_064_)
  );
  NAND _067_ (
    .A(\data1_i[21] ),
    .B(_063_),
    .Y(_000_)
  );
  NAND _068_ (
    .A(_064_),
    .B(_000_),
    .Y(\data_o[21] )
  );
  NAND _069_ (
    .A(select_i),
    .B(\data2_i[22] ),
    .Y(_001_)
  );
  NAND _070_ (
    .A(_063_),
    .B(\data1_i[22] ),
    .Y(_002_)
  );
  NAND _071_ (
    .A(_001_),
    .B(_002_),
    .Y(\data_o[22] )
  );
  NAND _072_ (
    .A(select_i),
    .B(\data2_i[23] ),
    .Y(_003_)
  );
  NAND _073_ (
    .A(_063_),
    .B(\data1_i[23] ),
    .Y(_004_)
  );
  NAND _074_ (
    .A(_003_),
    .B(_004_),
    .Y(\data_o[23] )
  );
  NAND _075_ (
    .A(select_i),
    .B(\data2_i[24] ),
    .Y(_005_)
  );
  NAND _076_ (
    .A(_063_),
    .B(\data1_i[24] ),
    .Y(_006_)
  );
  NAND _077_ (
    .A(_005_),
    .B(_006_),
    .Y(\data_o[24] )
  );
  NAND _078_ (
    .A(select_i),
    .B(\data2_i[25] ),
    .Y(_007_)
  );
  NAND _079_ (
    .A(_063_),
    .B(\data1_i[25] ),
    .Y(_008_)
  );
  NAND _080_ (
    .A(_007_),
    .B(_008_),
    .Y(\data_o[25] )
  );
  NAND _081_ (
    .A(select_i),
    .B(\data2_i[26] ),
    .Y(_009_)
  );
  NAND _082_ (
    .A(_063_),
    .B(\data1_i[26] ),
    .Y(_010_)
  );
  NAND _083_ (
    .A(_009_),
    .B(_010_),
    .Y(\data_o[26] )
  );
  NAND _084_ (
    .A(select_i),
    .B(\data2_i[27] ),
    .Y(_011_)
  );
  NAND _085_ (
    .A(_063_),
    .B(\data1_i[27] ),
    .Y(_012_)
  );
  NAND _086_ (
    .A(_011_),
    .B(_012_),
    .Y(\data_o[27] )
  );
  NAND _087_ (
    .A(select_i),
    .B(\data2_i[28] ),
    .Y(_013_)
  );
  NAND _088_ (
    .A(_063_),
    .B(\data1_i[28] ),
    .Y(_014_)
  );
  NAND _089_ (
    .A(_013_),
    .B(_014_),
    .Y(\data_o[28] )
  );
  NAND _090_ (
    .A(select_i),
    .B(\data2_i[29] ),
    .Y(_015_)
  );
  NAND _091_ (
    .A(_063_),
    .B(\data1_i[29] ),
    .Y(_016_)
  );
  NAND _092_ (
    .A(_015_),
    .B(_016_),
    .Y(\data_o[29] )
  );
  NAND _093_ (
    .A(select_i),
    .B(\data2_i[30] ),
    .Y(_017_)
  );
  NAND _094_ (
    .A(_063_),
    .B(\data1_i[30] ),
    .Y(_018_)
  );
  NAND _095_ (
    .A(_017_),
    .B(_018_),
    .Y(\data_o[30] )
  );
  NAND _096_ (
    .A(select_i),
    .B(\data2_i[31] ),
    .Y(_019_)
  );
  NAND _097_ (
    .A(_063_),
    .B(\data1_i[31] ),
    .Y(_020_)
  );
  NAND _098_ (
    .A(_019_),
    .B(_020_),
    .Y(\data_o[31] )
  );
  NAND _099_ (
    .A(select_i),
    .B(\data2_i[0] ),
    .Y(_021_)
  );
  NAND _100_ (
    .A(_063_),
    .B(\data1_i[0] ),
    .Y(_022_)
  );
  NAND _101_ (
    .A(_021_),
    .B(_022_),
    .Y(\data_o[0] )
  );
  NAND _102_ (
    .A(select_i),
    .B(\data2_i[1] ),
    .Y(_023_)
  );
  NAND _103_ (
    .A(_063_),
    .B(\data1_i[1] ),
    .Y(_024_)
  );
  NAND _104_ (
    .A(_023_),
    .B(_024_),
    .Y(\data_o[1] )
  );
  NAND _105_ (
    .A(select_i),
    .B(\data2_i[2] ),
    .Y(_025_)
  );
  NAND _106_ (
    .A(_063_),
    .B(\data1_i[2] ),
    .Y(_026_)
  );
  NAND _107_ (
    .A(_025_),
    .B(_026_),
    .Y(\data_o[2] )
  );
  NAND _108_ (
    .A(select_i),
    .B(\data2_i[3] ),
    .Y(_027_)
  );
  NAND _109_ (
    .A(_063_),
    .B(\data1_i[3] ),
    .Y(_028_)
  );
  NAND _110_ (
    .A(_027_),
    .B(_028_),
    .Y(\data_o[3] )
  );
  NAND _111_ (
    .A(select_i),
    .B(\data2_i[4] ),
    .Y(_029_)
  );
  NAND _112_ (
    .A(_063_),
    .B(\data1_i[4] ),
    .Y(_030_)
  );
  NAND _113_ (
    .A(_029_),
    .B(_030_),
    .Y(\data_o[4] )
  );
  NAND _114_ (
    .A(select_i),
    .B(\data2_i[5] ),
    .Y(_031_)
  );
  NAND _115_ (
    .A(_063_),
    .B(\data1_i[5] ),
    .Y(_032_)
  );
  NAND _116_ (
    .A(_031_),
    .B(_032_),
    .Y(\data_o[5] )
  );
  NAND _117_ (
    .A(select_i),
    .B(\data2_i[6] ),
    .Y(_033_)
  );
  NAND _118_ (
    .A(_063_),
    .B(\data1_i[6] ),
    .Y(_034_)
  );
  NAND _119_ (
    .A(_033_),
    .B(_034_),
    .Y(\data_o[6] )
  );
  NAND _120_ (
    .A(select_i),
    .B(\data2_i[7] ),
    .Y(_035_)
  );
  NAND _121_ (
    .A(_063_),
    .B(\data1_i[7] ),
    .Y(_036_)
  );
  NAND _122_ (
    .A(_035_),
    .B(_036_),
    .Y(\data_o[7] )
  );
  NAND _123_ (
    .A(select_i),
    .B(\data2_i[8] ),
    .Y(_037_)
  );
  NAND _124_ (
    .A(_063_),
    .B(\data1_i[8] ),
    .Y(_038_)
  );
  NAND _125_ (
    .A(_037_),
    .B(_038_),
    .Y(\data_o[8] )
  );
  NAND _126_ (
    .A(select_i),
    .B(\data2_i[9] ),
    .Y(_039_)
  );
  NAND _127_ (
    .A(_063_),
    .B(\data1_i[9] ),
    .Y(_040_)
  );
  NAND _128_ (
    .A(_039_),
    .B(_040_),
    .Y(\data_o[9] )
  );
  NAND _129_ (
    .A(select_i),
    .B(\data2_i[10] ),
    .Y(_041_)
  );
  NAND _130_ (
    .A(_063_),
    .B(\data1_i[10] ),
    .Y(_042_)
  );
  NAND _131_ (
    .A(_041_),
    .B(_042_),
    .Y(\data_o[10] )
  );
  NAND _132_ (
    .A(select_i),
    .B(\data2_i[11] ),
    .Y(_043_)
  );
  NAND _133_ (
    .A(_063_),
    .B(\data1_i[11] ),
    .Y(_044_)
  );
  NAND _134_ (
    .A(_043_),
    .B(_044_),
    .Y(\data_o[11] )
  );
  NAND _135_ (
    .A(select_i),
    .B(\data2_i[12] ),
    .Y(_045_)
  );
  NAND _136_ (
    .A(_063_),
    .B(\data1_i[12] ),
    .Y(_046_)
  );
  NAND _137_ (
    .A(_045_),
    .B(_046_),
    .Y(\data_o[12] )
  );
  NAND _138_ (
    .A(select_i),
    .B(\data2_i[13] ),
    .Y(_047_)
  );
  NAND _139_ (
    .A(_063_),
    .B(\data1_i[13] ),
    .Y(_048_)
  );
  NAND _140_ (
    .A(_047_),
    .B(_048_),
    .Y(\data_o[13] )
  );
  NAND _141_ (
    .A(select_i),
    .B(\data2_i[14] ),
    .Y(_049_)
  );
  NAND _142_ (
    .A(_063_),
    .B(\data1_i[14] ),
    .Y(_050_)
  );
  NAND _143_ (
    .A(_049_),
    .B(_050_),
    .Y(\data_o[14] )
  );
  NAND _144_ (
    .A(select_i),
    .B(\data2_i[15] ),
    .Y(_051_)
  );
  NAND _145_ (
    .A(_063_),
    .B(\data1_i[15] ),
    .Y(_052_)
  );
  NAND _146_ (
    .A(_051_),
    .B(_052_),
    .Y(\data_o[15] )
  );
  NAND _147_ (
    .A(select_i),
    .B(\data2_i[16] ),
    .Y(_053_)
  );
  NAND _148_ (
    .A(_063_),
    .B(\data1_i[16] ),
    .Y(_054_)
  );
  NAND _149_ (
    .A(_053_),
    .B(_054_),
    .Y(\data_o[16] )
  );
  NAND _150_ (
    .A(select_i),
    .B(\data2_i[17] ),
    .Y(_055_)
  );
  NAND _151_ (
    .A(_063_),
    .B(\data1_i[17] ),
    .Y(_056_)
  );
  NAND _152_ (
    .A(_055_),
    .B(_056_),
    .Y(\data_o[17] )
  );
  NAND _153_ (
    .A(select_i),
    .B(\data2_i[18] ),
    .Y(_057_)
  );
  NAND _154_ (
    .A(_063_),
    .B(\data1_i[18] ),
    .Y(_058_)
  );
  NAND _155_ (
    .A(_057_),
    .B(_058_),
    .Y(\data_o[18] )
  );
  NAND _156_ (
    .A(select_i),
    .B(\data2_i[19] ),
    .Y(_059_)
  );
  NAND _157_ (
    .A(_063_),
    .B(\data1_i[19] ),
    .Y(_060_)
  );
  NAND _158_ (
    .A(_059_),
    .B(_060_),
    .Y(\data_o[19] )
  );
  NAND _159_ (
    .A(select_i),
    .B(\data2_i[20] ),
    .Y(_061_)
  );
  NAND _160_ (
    .A(_063_),
    .B(\data1_i[20] ),
    .Y(_062_)
  );
  NAND _161_ (
    .A(_061_),
    .B(_062_),
    .Y(\data_o[20] )
  );
endmodule
